module top();
endmodule